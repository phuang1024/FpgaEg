module egcoding(
	input wire clk,
	input wire rst,
	input wire rx,
	input wire tx
);
endmodule